module insertionSort #(
    parameter NUM_VALS = 5,
    parameter SIZE_DATA = 8
)(
    input  logic                         i_clk,
    input  logic                         i_rst_n,
    input  logic                         i_start,
    input  logic [NUM_VALS*SIZE_DATA-1:0] i_data,
    output logic                         o_done,
    output logic [NUM_VALS*SIZE_DATA-1:0] o_data
);

    // State encoding
    typedef enum logic [2:0] {
        b0, // Reset/init
        b1, // Load data into internal array
        b2, // Wait for start
        b3, // Use compare_block for first two elements
        b4, // Select key
        b5, // While loop condition
        b6, // Shift and insert
        b7  // Done
    } state_t;

    state_t state;

    // Internal array
    logic [SIZE_DATA-1:0] arr_temp [NUM_VALS-1:0];
    logic [SIZE_DATA-1:0] key;
    int i_sign; // current index of insertion

    // Compare block outputs
    logic [SIZE_DATA-1:0] w_less_data;
    logic [SIZE_DATA-1:0] w_greater_data;

    // FSM & datapath
    always_ff @(posedge i_clk or negedge i_rst_n) begin
        if (!i_rst_n) begin
            state <= b0;
            o_done <= 1'b0;
            i_sign <= 0;
        end else begin
            case (state)
                b0: begin
                    o_done <= 1'b0;
                    state <= b1;
                end

                b1: begin
                    // Load input data to internal array
                    for (int i = 0; i < NUM_VALS; i++) begin
                        arr_temp[i] <= i_data[i*SIZE_DATA +: SIZE_DATA];
                    end
                    state <= b2;
                end

                b2: begin
                    // Wait for start signal
                    if (i_start)
                        state <= b3;
                end

                b3: begin
                    // Use compare_block to sort first 2 elements
                    arr_temp[0] <= w_less_data;
                    arr_temp[1] <= w_greater_data;
                    i_sign <= 2; // Start insertion from 3rd element
                    state <= b4;
                end

                b4: begin
                    if (i_sign < NUM_VALS) begin
                        key <= arr_temp[i_sign];
                        i_sign <= i_sign - 1;
                        state <= b5;
                    end else begin
                        state <= b7;
                    end
                end

                b5: begin
                    if ((i_sign >= 0) && (key < arr_temp[i_sign])) begin
                        arr_temp[i_sign + 1] <= arr_temp[i_sign];
                        i_sign <= i_sign - 1;
                        state <= b5; // Repeat
                    end else begin
                        state <= b6;
                    end
                end

                b6: begin
                    arr_temp[i_sign + 1] <= key;
                    i_sign <= i_sign + 2;
                    state <= b4;
                end

                b7: begin
                    // Sorting done
                    for (int i = 0; i < NUM_VALS; i++) begin
                        o_data[i*SIZE_DATA +: SIZE_DATA] <= arr_temp[i];
                    end
                    o_done <= 1'b1;
                    state <= b0; // reset for next run
                end

                default: state <= b0;
            endcase
        end
    end

    // === Compare block instantiation ===
    compare_block #(
        .SIZE_DATA(SIZE_DATA)
    ) u_compare_block (
        .i_data_a(arr_temp[0]),
        .i_data_b(arr_temp[1]),
        .i_mode(1'b0),
        .o_less_data(w_less_data),
        .o_greater_data(w_greater_data)
    );

endmodule

// module insertionSort #(
//     parameter SIZE_DATA = 8,
//     parameter NUM_VALS  = 8
// )(
//     input  logic                     i_clk       ,
//     input  logic                     i_rst_n     ,
//     input  logic                     i_start     ,
//     input  logic                     i_mode      , // 0: ascending, 1: descending 
    // input  logic [SIZE_DATA-1:0]     i_data [NUM_VALS],
    // output logic [SIZE_DATA-1:0]     o_data [NUM_VALS],
//     output logic                     o_done
// );

// logic [SIZE_DATA-1:0] arr_temp [NUM_VALS];
// logic [SIZE_DATA-1:0] w_temp_data_0, w_temp_data_1;

// compare_block #(
//     .SIZE_DATA(SIZE_DATA)
// ) u_compare_block (
//     .i_data_a(i_data[0]),
//     .i_data_b(i_data[1]),
//     .i_mode(i_mode),
//     .o_less_data(w_temp_data_0),
//     .o_greater_data(w_temp_data_1)
// );

// always_ff @(posedge i_clk or negedge i_rst_n) begin : proc_two_ele_first
//     if(~i_rst_n) begin
//         for(int i = 0; i < NUM_VALS; i ++) begin
//             arr_temp[i] <= '0;
//         end
//     end else if(state == LOAD_I) begin
//         arr_temp[0] <= w_temp_data_0;
//         arr_temp[1] <= w_temp_data_1;
//         for(int i = 2; i < NUM_VALS; i ++) begin
//             arr_temp[i] <= i_data[i];
//         end
//     end else if(state == LOAD_J) begin
//         arr_temp[j_sign + 1'b1] <= arr_temp[j_sign];
//     end else if(state == INSERT) begin
//         arr_temp[j_sign + 1'b1] <= key;
//     end
// end

// typedef enum logic [2:0] { 
//     IDLE        ,
//     LOAD_I      ,
//     COMPARE_I   ,
//     LOAD_J      ,
//     COMPARE_J   ,
//     INSERT      ,
//     DONE        
// } state_t;

// state_t state, n_state;

// logic [$clog2(SIZE_DATA)-1:0] i_sign;
// logic [$clog2(NUM_VALS)-1:0] j_sign;
// logic [SIZE_DATA-1:0] key;

// logic w_update_compare_i, w_update_load_j;
// assign w_update_compare_i = (i_sign < NUM_VALS);
// assign w_update_load_j = (i_mode) ? (key > arr_temp[j_sign]) : (key < arr_temp[j_sign]);

// always_comb begin : proc_next_state
//     case(state)
//         IDLE:        n_state = (i_start) ? LOAD_I : IDLE;
//         LOAD_I:      n_state = COMPARE_I;
//         COMPARE_I:   n_state = (w_update_compare_i) ? LOAD_J : DONE;
//         LOAD_J:      n_state = (j_sign != 0 && w_update_load_j) ? COMPARE_J : INSERT;
//         COMPARE_J:   n_state = LOAD_J;
//         INSERT:      n_state = COMPARE_I;
//         DONE:        n_state = IDLE;
//         default:     n_state = IDLE;
//     endcase
// end

// always_ff @(posedge i_clk or negedge i_rst_n) begin
//     if(~i_rst_n) begin
//         i_sign <= 2;
//         j_sign <= '0;
//         key    <= '0;
//         o_done <= '0;
//         state  <= IDLE;
//     end else begin
//         state <= n_state;
//         case(state)
//             IDLE: begin
//                 i_sign <= 2;
//                 j_sign <= '0;
//                 key    <= '0;
//                 o_done <= '0;
//             end
//             LOAD_I: begin
//                 i_sign <= 2;
//                 j_sign <= '0;
//                 key    <= '0;
//                 o_done <= '0;
//             end
//             COMPARE_I: begin
//                 j_sign <= i_sign - 1'b1;
//                 key    <= arr_temp[i_sign];
//             end
//             COMPARE_J: begin
//                 j_sign <= j_sign - 1'b1;
//             end
//             INSERT: begin
//                 i_sign <= i_sign + 1'b1;
//             end
//             DONE: begin
//                 i_sign <= 2;
//                 j_sign <= '0;
//                 key    <= '0;
//                 o_done <= 1'b1;
//             end
//             default: begin
//                 o_done <= 1'b0;
//             end
//         endcase
//     end
// end

// always_ff @(posedge i_clk or negedge i_rst_n) begin
//     if(~i_rst_n) begin
//         for(int i = 0; i < NUM_VALS; i++) begin
//             o_data[i] <= '0;
//         end
//     end else if(o_done) begin
//         for(int i = 0; i < NUM_VALS; i++) begin
//             o_data[i] <= arr_temp[i];
//         end
//     end
// end

// endmodule
// module insertionSort #(
//     parameter NUM_VALS = 5,
//     parameter SIZE_DATA = 8
// )(
//     input  logic                         i_clk,
//     input  logic                         i_rst_n,
//     input  logic                         i_start,
//     input  logic [SIZE_DATA-1:0]         i_data [NUM_VALS],
//     output logic                         o_done,
//     output logic [SIZE_DATA-1:0]         o_data [NUM_VALS]
// );

//     // State encoding
//     typedef enum logic [2:0] {
//         b0, // Reset/init
//         b1, // Load data into internal array
//         b2, // Wait for start
//         b3, // Use compare_block for first two elements
//         b4, // Select key
//         b5, // While loop condition
//         b6, // Shift and insert
//         b7  // Done
//     } state_t;

//     state_t state;

//     // Internal array
//     logic [SIZE_DATA-1:0] arr_temp [NUM_VALS];
//     logic [SIZE_DATA-1:0] key;
//     int i_sign;

//     // Compare block outputs
//     logic [SIZE_DATA-1:0] w_less_data;
//     logic [SIZE_DATA-1:0] w_greater_data;

//     // FSM & datapath
//     always_ff @(posedge i_clk or negedge i_rst_n) begin
//         if (!i_rst_n) begin
//             state   <= b0;
//             o_done  <= 1'b0;
//             i_sign  <= 0;
//         end else begin
//             case (state)
//                 b0: begin
//                     o_done <= 1'b0;
//                     state  <= b1;
//                 end

//                 b1: begin
//                     // Load input data to internal array
//                     for (int i = 0; i < NUM_VALS; i++) begin
//                         arr_temp[i] <= i_data[i];
//                     end
//                     state <= b2;
//                 end

//                 b2: begin
//                     // Wait for start signal
//                     if (i_start)
//                         state <= b3;
//                 end

//                 b3: begin
//                     // Use compare_block to sort first 2 elements
//                     arr_temp[0] <= w_less_data;
//                     arr_temp[1] <= w_greater_data;
//                     i_sign      <= 2;
//                     state       <= b4;
//                 end

//                 b4: begin
//                     if (i_sign < NUM_VALS) begin
//                         key    <= arr_temp[i_sign];
//                         i_sign <= i_sign - 1;
//                         state  <= b5;
//                     end else begin
//                         state <= b7;
//                     end
//                 end

//                 b5: begin
//                     if ((i_sign >= 0) && (key < arr_temp[i_sign])) begin
//                         arr_temp[i_sign + 1] <= arr_temp[i_sign];
//                         i_sign <= i_sign - 1;
//                         state  <= b5;
//                     end else begin
//                         state <= b6;
//                     end
//                 end

//                 b6: begin
//                     arr_temp[i_sign + 1] <= key;
//                     i_sign <= i_sign + 2;
//                     state  <= b4;
//                 end

//                 b7: begin
//                     for (int i = 0; i < NUM_VALS; i++) begin
//                         o_data[i] <= arr_temp[i];
//                     end
//                     o_done <= 1'b1;
//                     state  <= b0;
//                 end

//                 default: state <= b0;
//             endcase
//         end
//     end

//     // === Compare block instantiation ===
//     compare_block #(
//         .SIZE_DATA(SIZE_DATA)
//     ) u_compare_block (
//         .i_data_a(arr_temp[0]),
//         .i_data_b(arr_temp[1]),
//         .i_mode(1'b0), // ascending
//         .o_less_data(w_less_data),
//         .o_greater_data(w_greater_data)
//     );

// endmodule
