module PA_buf_greater #()();

endmodule
