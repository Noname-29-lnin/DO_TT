module Top_module(
    input logic                 i_clk       ,
    input logic                 i_rst_n     ,
    input logic                 i_start     ,
);

endmodule
