module PA_cal_depth_addr #(

)(

);

endmodule
