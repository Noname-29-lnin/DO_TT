module PA_partition #()();

endmodule
