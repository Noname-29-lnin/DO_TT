module DI_control #()();

endmodule
